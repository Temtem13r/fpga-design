`include "cpu.v"

module cpu_tb;

	initial begin
		
	end

endmodule